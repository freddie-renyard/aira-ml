parameter PRE_NEURON_NUM = <pre_neurons>,
POST_NEURON_NUM = <post_neurons>,

N_MAN_INPUT = <n_man_input>,
N_EXP_INPUT = <n_exp_input>,

N_MAN_WEIGHT = <n_man_weight>,
N_EXP_WEIGHT = <n_exp_weight>,

N_MAN_OUT = <n_man_out>,
N_EXP_OUT = <n_exp_out>,
    
N_OVERFLOW = <n_overflow>,
MULT_EXTRA = <mult_extra>,

MEM_DEPTH = <mem_depth>,
N_ADDR_DELTA = <n_delta>,

ACT_FUNC = <act_code>,

FILE_ID = <index>;
