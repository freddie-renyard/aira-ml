

    // Connection from object <i_pre> to top file output port 
    assign o_data = o_data_<i_pre>;
    assign o_d_valid = o_d_valid_<i_pre>;
    assign i_stall_<i_pre> = i_stall;