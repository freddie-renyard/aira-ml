// Layer <i> Common Parameters 
parameter N_MAN_INPUT_<i> = <n_man_input>,
N_EXP_INPUT_<i> = <n_exp_input>,
N_INPUT_<i> = <n_input>,

N_MAN_WEIGHT_<i> = <n_man_weight>,
N_EXP_WEIGHT_<i> = <n_exp_weight>,

N_MAN_OUT_<i> = <n_man_out>,
N_EXP_OUT_<i> = <n_exp_out>,
N_OUTPUT_<i> = <n_output>,
    
N_OVERFLOW_<i> = <n_overflow>,
MULT_EXTRA_<i> = <mult_extra>;

