// Module Input and Output parameters
parameter N_MODULE_INPUT = <n_mod_in>,
N_MODULE_OUTPUT = <n_mod_out>;

