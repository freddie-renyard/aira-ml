parameter PRE_NEURON_NUM_<i> = <pre_neurons>,
POST_NEURON_NUM_<i> = <post_neurons>,

N_MAN_INPUT_<i> = <n_man_input>,
N_EXP_INPUT_<i> = <n_exp_input>,

N_MAN_WEIGHT_<i> = <n_man_weight>,
N_EXP_WEIGHT_<i> = <n_exp_weight>,

N_MAN_OUT_<i> = <n_man_out>,
N_EXP_OUT_<i> = <n_exp_out>,
    
N_OVERFLOW_<i> = <n_overflow>,
MULT_EXTRA_<i> = <mult_extra>,

MEM_DEPTH_<i> = <mem_depth>,
N_ADDR_DELTA_<i> = <n_delta>,

ACT_FUNC_<i> = <act_code>,

FILE_ID_<i> = <i>;
