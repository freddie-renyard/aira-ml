    
    
    // Dense Layer <i> Wires
    wire [N_INPUT_<i>-1:0] i_data_<i>;
    wire i_d_valid_<i>;
    wire o_stall_<i>;
    
    wire [N_OUTPUT_<i>-1:0] o_data_<i>;
    wire o_d_valid_<i>;
    wire i_stall_<i>;